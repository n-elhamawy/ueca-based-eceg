/*Elliptic Curve parameters y^2 = x^2 + Ax + B
  modulo the prime p
  with the bit length DATAWIDTH */

`define faultWidth  8
 /*Parameters for Elliptic Curve with 521 bits*/

`define DATAWIDTH  521
`define p          521'd6864797660130609714981900799081393217269435300143305409394463459185543183397656052122559640661454554977296311391480858037121987999716643812574028291115057151
`define A          521'd6864797660130609714981900799081393217269435300143305409394463459185543183397656052122559640661454554977296311391480858037121987999716643812574028291115057148
`define B          521'd1093849038073734274511112390766805569936207598951683748994586394495953116150735016013708737573759623248592132296706313309438452531591012912142327488478985984
`define Px         521'd2661740802050217063228768716723360960729859168756973147706671368418802944996427808491545080627771902352094241225065558662157113545570916814161637315895999846
`define Py         521'd3757180025770020463545507224491183603594455134769762486694567779615544477440556316691234405012945539562144444537289428522585666729196580810124344277578376784
`define Mx0        521'd6581699809797034456215217677504225167184642460997740611822024977354528670332877711961660616359114018821487277280083055191025738601442093308170769130244837783
`define My0        521'd1997278802466087953174121891499340641274644866423460163424047421289940218188598764635249404031736012724075294139346145992226211508304690854187362956785301376
`define secretKey  521'd171721461964413649154124237231217104981741483823050811371748171477717014312117918713257571422061672202172011381723911493166641091712291841619622916424923524 
`define k          521'd591851771144408419225413818146254719913217193917790199118713275178137521610413522142549722247641591351802421144551918596120198176101722551951252461273690240

 /*Parameters for Elliptic Curve with 384 bits*/
 /*
`define DATAWIDTH  384
`define p          384'd39402006196394479212279040100143613805079739270465446667948293404245721771496870329047266088258938001861606973112319
`define A          384'd39402006196394479212279040100143613805079739270465446667948293404245721771496870329047266088258938001861606973112316
`define B          384'd27580193559959705877849011840389048093056905856361568521428707301988689241309860865136260764883745107765439761230575
`define Px         384'd26247035095799689268623156744566981891852923491109213387815615900925518854738050089022388053975719786650872476732087
`define Py         384'd8325710961489029985546751289520108179287853048861315594709205902480503199884419224438643760392947333078086511627871
`define Mx0        384'd5273320726046279714052782309791752925190860505809940144458899488645531928156241880041348929390131490907893417210083
`define My0        384'd26655923019261778224161832290008317559844283029247519399262162425172313950821409655533332657708521002737382803200618
`define secretKey  384'd1151194113898485231351361931212372924716043197771792051507014026175212232252371963158127121562020316321319013287260
`define k          384'd2343731562532222193168217122615838024018598107101811568316015818734159164412162229131218129223186321773312219104112 
*/

    /*Parameters for Elliptic Curve with 256 bits*/
/*
`define DATAWIDTH  256
`define p          256'd115792089210356248762697446949407573530086143415290314195533631308867097853951
`define A          256'd115792089210356248762697446949407573530086143415290314195533631308867097853948
`define B          256'd41058363725152142129326129780047268409114441015993725554835256314039467401291
`define Px         256'd48439561293906451759052585252797914202762949526041747995844080717082404635286
`define Py         256'd36134250956749795798585127919587881956611106672985015071877198253568414405109
`define Mx0        256'd72649262508960331895015918013687691681933102559554532061209154701483247778628
`define My0        256'd88449348244875801639180290383169546753923522234842718834683349047530142861915
`define secretKey  256'd302296273192362411826411822524524874196150110112821521380941085611523125149 
`define k          256'd772261881201649925251206127625024610416622894731981201117353782358518219152 

*/

   /*Parameters for Elliptic Curve with 224 bits*/
/*
`define DATAWIDTH  224
`define p          224'd26959946667150639794667015087019630673557916260026308143510066298881
`define A          224'd26959946667150639794667015087019630673557916260026308143510066298878
`define B          224'd18958286285566608000408668544493926415504680968679321075787234672564
`define Px         224'd19277929113566293071110308034699488026831934219452440156649784352033
`define Py         224'd19926808758034470970197974289220981123180760759394043754012972449332
`define Mx0        224'd26544976231971333689576543919985296373708387637830311523141116612874
`define My0        224'd8364236922062653245278732495200776517634578356291150317373038179662
`define secretKey  224'd355623414112510197227313258115522153242124190217172561511411019020
`define k          224'd12315014760664494110118213157591421782231625418617247910714524520210 
 */
  /*Parameters for Elliptic Curve with 192 bits*/
/*
`define DATAWIDTH  192
`define p          192'd6277101735386680763835789423207666416083908700390324961279
`define A          192'd6277101735386680763835789423207666416083908700390324961276
`define B          192'd2455155546008943817740293915197451784769108058161191238065
`define Px         192'd602046282375688656758213480587526111916698976636884684818
`define Py         192'd174050332293622031404857552280219410364023488927386650641
`define Mx0        192'd605531991447545055930502119775989644341093705383285943229
`define My0        192'd5390682307141156010169044267689660431108249307394684532795
`define secretKey  192'd2063415921261422524613818319217472531059261595414616152 
`define k          192'd1337425231106111949616166212841322013811222231098185242 
 */
 /*Parameters for Elliptic Curve with 160 bits*/
/*
`define DATAWIDTH  160
`define p          160'd1461501637330902918203684832716283019653785059327
`define A          160'd1461501637330902918203684832716283019653785059324
`define B          160'd163235791306168110546604919403271579530548345413
`define Px         160'd425826231723888350446541592701409065913635568770
`define Py         160'd203520114162904107873991457957346892027982641970
`define Mx0        160'd622767356176297183435784449477825205923203789449
`define My0        160'd132078438334177474887606962011735303624788231865
`define secretKey  160'd154143153762283812959131661311816348581221164337 
`define k          160'd148489441658014101902542261612178131771619314440 
*/

/*Parameters for Elliptic Curve with 128 bits*/
/*
`define DATAWIDTH  128
`define p          128'd340282366762482138434845932244680310783
`define A          128'd340282366762482138434845932244680310780
`define B          128'd308990863222245658030922601041482374867
`define Px         128'd29408993404948928992877151431649155974
`define Py         128'd275621562871047521857442314737465260675
`define Mx0        128'd25022131429364248112951584293624460930
`define My0        128'd121817100096969938286892229223484993851
`define secretKey  128'd42624822515914917023322916317892122324 
//`define secretKey  128'd2075174161569616921896229281511211628  
`define k          128'd166841011151241872031651641266734614613           
*/

/*Parameters for Elliptic Curve with 15 bits*/
/*
`define DATAWIDTH   15
`define p           15'd32003
`define A           15'd18786
`define B           15'd12857
`define Px          15'd16533
`define Py          15'd31897
`define Mx0         15'd16775
`define My0         15'd20887
`define secretKey   15'd23413
`define k           15'd15321
*/
